module pwm(

);

endmodule